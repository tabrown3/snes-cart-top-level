module cmd_manager
(
    input clk,
    input [7:0] in_byte,
    input byte_finished
);

endmodule