module cmd_manager
(
    input clk,
    input [7:0] in_byte,
    input byte_finished,
    output [7:0] out_byte = 8'h00
);

endmodule